
//# sourceMappingURL=async_fifo_reset_sync.sv.map
