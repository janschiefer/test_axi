///AXI4 bus package prototype









//# sourceMappingURL=axi_if.sv.map
