

//# sourceMappingURL=async_fifo.sv.map
