
/// Asynchronous handshake
///
/// Asynchronous data transmitter based on handshake protocol.
/// Generic parameter `S` is a module name of synchrinoizer.

//# sourceMappingURL=async_handshake.sv.map
