
//# sourceMappingURL=synchronizer.sv.map
